---------------------------------------------------------------------------------
--
-- Copyright (c) 2017 by VLSI Systems Design Laboratory,
-- The University of Engineering and Technology, Vietnam National University.
-- All right resevered.
--
-- Copyright notification
-- No part may be reproduced except as authorized by written permission.
-- 
-- @File            : NN_selector.vhd
-- @Author          : Xuan-Thuan Nguyen 	 @Modifier           :
-- @Created Date    :   /  /      		 @Modified Date      :
-- @Project         : Library
-- @Module          : NN_selector
-- @Description     : Description of module.
-- @Version         : 0.1beta
-- @ID              : N/A
--
--------------------------------------------------------------------------------

---------------------------------------------------------------------------------
-- Library declaration
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
---------------------------------------------------------------------------------
-- Entity declaration
--------------------------------------------------------------------------------- 
entity selecctor is
port
(
	clk 			: in 	std_logic;  
	areset 			: in 	std_logic;  
	enable_update 	: out 	std_logic  
);
end selecctor; 

---------------------------------------------------------------------------------
-- Architecture description
---------------------------------------------------------------------------------
architecture beh of selecctor is
constant N : integer :=13;
signal counter : signed(7 downto 0);
begin
	count :process(clk, areset)
			begin
				if(rising_edge(clk)) then
					if(areset = '1') then
						counter <= (others => '0');
					else
						if(counter = to_signed((N-1),8)) then
							counter <= (others => '0');
						else
							counter <= counter + to_signed(1,8);
						end if;
					end if;
				end if;
			end process count;
	enb_upd:process(clk, areset)
			begin
				if(rising_edge(clk)) then
					if(areset = '1') then
						enable_update <= '0';
					else
						if(counter = to_signed((N-1),8)) then
							enable_update <= '1';
						else
							enable_update <= '0';
						end if;
					end if;
				end if;
			end process enb_upd;
end beh;
