`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:37:14 10/13/2017
// Design Name:   backward
// Module Name:   C:/Users/igarashi/Desktop/20171013_1442_backward/backward/backward_tb.v
// Project Name:  backward
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: backward
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module backward_tb;

	// Inputs
	reg clk;
	reg res;
	reg [31:0] a3_1;
	reg [31:0] a3_2;
	reg [31:0] a2_1;
	reg [31:0] a2_2;
	reg [31:0] a2_3;
	reg [31:0] k_1;
	reg [31:0] k_2;
	reg [31:0] t_1;
	reg [31:0] t_2;
	reg [31:0] w3_11;
	reg [31:0] w3_21;
	reg [31:0] w3_31;
	reg [31:0] w3_12;
	reg [31:0] w3_22;
	reg [31:0] w3_32;

	// Outputs
	wire [31:0] cap_delta_w3_11;
	wire [31:0] cap_delta_w3_21;
	wire [31:0] cap_delta_w3_31;
	wire [31:0] cap_delta_w3_12;
	wire [31:0] cap_delta_w3_22;
	wire [31:0] cap_delta_w3_32;
	wire [31:0] cap_delta_w2_11;
	wire [31:0] cap_delta_w2_21;
	wire [31:0] cap_delta_w2_12;
	wire [31:0] cap_delta_w2_22;
	wire [31:0] cap_delta_w2_13;
	wire [31:0] cap_delta_w2_23;
	wire [31:0] cap_delta_b3_1;
	wire [31:0] cap_delta_b3_2;
	wire [31:0] cap_delta_b2_1;
	wire [31:0] cap_delta_b2_2;
	wire [31:0] cap_delta_b2_3;

	// Instantiate the Unit Under Test (UUT)
	backward uut (
		.clk(clk), 
		.res(res), 
		.a3_1(a3_1), 
		.a3_2(a3_2), 
		.a2_1(a2_1), 
		.a2_2(a2_2), 
		.a2_3(a2_3), 
		.k_1(k_1), 
		.k_2(k_2), 
		.t_1(t_1), 
		.t_2(t_2), 
		.w3_11(w3_11), 
		.w3_21(w3_21), 
		.w3_31(w3_31), 
		.w3_12(w3_12), 
		.w3_22(w3_22), 
		.w3_32(w3_32), 
		.cap_delta_w3_11(cap_delta_w3_11), 
		.cap_delta_w3_21(cap_delta_w3_21), 
		.cap_delta_w3_31(cap_delta_w3_31), 
		.cap_delta_w3_12(cap_delta_w3_12), 
		.cap_delta_w3_22(cap_delta_w3_22), 
		.cap_delta_w3_32(cap_delta_w3_32), 
		.cap_delta_w2_11(cap_delta_w2_11), 
		.cap_delta_w2_21(cap_delta_w2_21), 
		.cap_delta_w2_12(cap_delta_w2_12), 
		.cap_delta_w2_22(cap_delta_w2_22), 
		.cap_delta_w2_13(cap_delta_w2_13), 
		.cap_delta_w2_23(cap_delta_w2_23), 
		.cap_delta_b3_1(cap_delta_b3_1), 
		.cap_delta_b3_2(cap_delta_b3_2), 
		.cap_delta_b2_1(cap_delta_b2_1), 
		.cap_delta_b2_2(cap_delta_b2_2), 
		.cap_delta_b2_3(cap_delta_b2_3)
	);

	parameter STEP = 100;
	
	always begin
		clk = 1; #(STEP/2);
		clk = 0; #(STEP/2);
	end


	initial begin
		// Initialize Inputs
		res = 0;
		a3_1 = 0;
		a3_2 = 0;
		a2_1 = 0;
		a2_2 = 0;
		a2_3 = 0;
		k_1 = 0;
		k_2 = 0;
		t_1 = 0;
		t_2 = 0;
		w3_11 = 0;
		w3_21 = 0;
		w3_31 = 0;
		w3_12 = 0;
		w3_22 = 0;
		w3_32 = 0;

		#50
		res = 1;
		#STEP
		res = 0;
		//#(STEP*20)
		//(8,8)
		#(STEP*10) 
		a3_1 	= 32'b0000_0000_1111_1110_0010_1101_0100_1010; 
		a3_2 	= 32'b0000_0000_1111_1101_1010_1001_1111_0001;
		a2_1 	= 32'b0000_0000_1111_1011_0001_1010_1011_0000;
		a2_2 	= 32'b0000_0000_1111_1111_1001_0000_1000_1011;
		a2_3 	= 32'b0000_0000_1111_1111_0000_0101_0101_1100;
		k_1   	= 32'b0000_1000_0000_0000_0000_0000_0000_0000; 
		k_2   	= 32'b0000_1000_0000_0000_0000_0000_0000_0000;
		t_1  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		w3_11 = 32'b0000_0000_0001_1001_1110_0001_1011_0010;
		w3_21 = 32'b0000_0000_0011_0011_0011_0011_0011_0011;
		w3_31 = 32'b0000_0001_0100_1100_1100_1100_1100_1100;
		w3_12 = 32'b0000_0000_0011_0011_0011_0011_0011_0011;
		w3_22 = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
		w3_32 = 32'b0000_0001_0001_1001_1001_1001_1001_1001;
		
		//(8,5)
		#STEP 
		a3_1 = 32'b00000000111010110110110110110001;
		a3_2 = 32'b00000000000000001100111111101101;
		a2_1 = 32'b00000000111100001001111000101001;
		a2_2 = 32'b00000000111111100000111101101011;
		a2_3 = 32'b00000000111111101010100111100101;
		k_1   = 32'b00001000000000000000000000000000;
		k_2   = 32'b00000101000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;

		//(5,8)
		#STEP 
		a3_1 = 32'b00000000111111111110001111001000;
		a3_2 = 32'b00000000111111010000001000010000;
		a2_1 = 32'b00000000111110011011111101101001;
		a2_2 = 32'b00000000111111101110010000100001;
		a2_3 = 32'b00000000111110100001111000101000;
		k_1   = 32'b00000101000000000000000000000000;
		k_2   = 32'b00001000000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		
		//(5,5)
		#STEP 
		a3_1 = 32'b00000000111111111101100101110000;
		a3_2 = 32'b00000000111100100101010000101001;
		a2_1 = 32'b00000000111010110110110110110001;
		a2_2 = 32'b00000000111110110001101010110000;
		a2_3 = 32'b00000000111110000000011011110101;
		k_1   = 32'b00000101000000000000000000000000;
		k_2   = 32'b00000101000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		
		#(STEP*10);

		//(8,8)
		#STEP 
		a3_1 	= 32'b0000_0000_1111_1110_0010_1101_0100_1010; 
		a3_2 	= 32'b0000_0000_1111_1101_1010_1001_1111_0001;
		a2_1 	= 32'b0000_0000_1111_1011_0001_1010_1011_0000;
		a2_2 	= 32'b0000_0000_1111_1111_1001_0000_1000_1011;
		a2_3 	= 32'b0000_0000_1111_1111_0000_0101_0101_1100;
		k_1   	= 32'b0000_1000_0000_0000_0000_0000_0000_0000; 
		k_2   	= 32'b0000_1000_0000_0000_0000_0000_0000_0000;
		t_1  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		w3_11 = 32'b0000_0000_0001_1001_1110_0001_1011_0010;
		w3_21 = 32'b0000_0000_0011_0011_0011_0011_0011_0011;
		w3_31 = 32'b0000_0001_0100_1100_1100_1100_1100_1100;
		w3_12 = 32'b0000_0000_0011_0011_0011_0011_0011_0011;
		w3_22 = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
		w3_32 = 32'b0000_0001_0001_1001_1001_1001_1001_1001;
		
		//(8,5)
		#STEP 
		a3_1 = 32'b00000000111010110110110110110001;
		a3_2 = 32'b00000000000000001100111111101101;
		a2_1 = 32'b00000000111100001001111000101001;
		a2_2 = 32'b00000000111111100000111101101011;
		a2_3 = 32'b00000000111111101010100111100101;
		k_1   = 32'b00001000000000000000000000000000;
		k_2   = 32'b00000101000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;

		//(5,8)
		#STEP 
		a3_1 = 32'b00000000111111111110001111001000;
		a3_2 = 32'b00000000111111010000001000010000;
		a2_1 = 32'b00000000111110011011111101101001;
		a2_2 = 32'b00000000111111101110010000100001;
		a2_3 = 32'b00000000111110100001111000101000;
		k_1   = 32'b00000101000000000000000000000000;
		k_2   = 32'b00001000000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		
		//(5,5)
		#STEP 
		a3_1 = 32'b00000000111111111101100101110000;
		a3_2 = 32'b00000000111100100101010000101001;
		a2_1 = 32'b00000000111010110110110110110001;
		a2_2 = 32'b00000000111110110001101010110000;
		a2_3 = 32'b00000000111110000000011011110101;
		k_1   = 32'b00000101000000000000000000000000;
		k_2   = 32'b00000101000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		
		#(STEP*10);

		//(8,8)
		#STEP 
		a3_1 	= 32'b0000_0000_1111_1110_0010_1101_0100_1010; 
		a3_2 	= 32'b0000_0000_1111_1101_1010_1001_1111_0001;
		a2_1 	= 32'b0000_0000_1111_1011_0001_1010_1011_0000;
		a2_2 	= 32'b0000_0000_1111_1111_1001_0000_1000_1011;
		a2_3 	= 32'b0000_0000_1111_1111_0000_0101_0101_1100;
		k_1   	= 32'b0000_1000_0000_0000_0000_0000_0000_0000; 
		k_2   	= 32'b0000_1000_0000_0000_0000_0000_0000_0000;
		t_1  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		w3_11 = 32'b0000_0000_0001_1001_1110_0001_1011_0010;
		w3_21 = 32'b0000_0000_0011_0011_0011_0011_0011_0011;
		w3_31 = 32'b0000_0001_0100_1100_1100_1100_1100_1100;
		w3_12 = 32'b0000_0000_0011_0011_0011_0011_0011_0011;
		w3_22 = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
		w3_32 = 32'b0000_0001_0001_1001_1001_1001_1001_1001;
		
		//(8,5)
		#STEP 
		a3_1 = 32'b00000000111010110110110110110001;
		a3_2 = 32'b00000000000000001100111111101101;
		a2_1 = 32'b00000000111100001001111000101001;
		a2_2 = 32'b00000000111111100000111101101011;
		a2_3 = 32'b00000000111111101010100111100101;
		k_1   = 32'b00001000000000000000000000000000;
		k_2   = 32'b00000101000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;

		//(5,8)
		#STEP 
		a3_1 = 32'b00000000111111111110001111001000;
		a3_2 = 32'b00000000111111010000001000010000;
		a2_1 = 32'b00000000111110011011111101101001;
		a2_2 = 32'b00000000111111101110010000100001;
		a2_3 = 32'b00000000111110100001111000101000;
		k_1   = 32'b00000101000000000000000000000000;
		k_2   = 32'b00001000000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		
		//(5,5)
		#STEP 
		a3_1 = 32'b00000000111111111101100101110000;
		a3_2 = 32'b00000000111100100101010000101001;
		a2_1 = 32'b00000000111010110110110110110001;
		a2_2 = 32'b00000000111110110001101010110000;
		a2_3 = 32'b00000000111110000000011011110101;
		k_1   = 32'b00000101000000000000000000000000;
		k_2   = 32'b00000101000000000000000000000000;
		t_1  	= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
		t_2  	= 32'b0000_0001_0000_0000_0000_0000_0000_0000;
		
		
		// Add stimulus here
	// End
	#(STEP*10) $finish;
	end
	endmodule


