`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Kyushu Institute of Technology
// Engineer: DSP Lab
// 
// Create Date:    13:48:25 09/06/2017 
// Design Name:    Neural Network (using backpropagation)
// Module Name:    mem
// Project Name:   LSI Design Contest in Okinawa 2018
// Target Devices: 
// Tool versions: 
//
// Description: 
// 	    8 bits memory to store value of sigmoid calculation
// Input:
//		clk	    : 1 bit
//		din 	: 1 bit : read enable
//		addr    : 8 bits 0000.0000 unsigned : value of sigmoid func with input from -8.0 to 7.93750 
// Output: 
//		dout	: 16 bits 00_0000.0000_0000_00 unsigned : output value for sigmoid func.
// Latency: 1 clk
// 
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Name : date : what changed
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mem(clk, din, addr, dout);
 parameter DWIDTH=16;								//bit width of data
 parameter AWIDTH=8;								//bit width of address
 parameter DWIDTH_TMP=32;
 
 input clk, din;									//	din : read enable signal
 input [AWIDTH-1:0] addr;							// 8 bits address [7:0]	addr
 output [DWIDTH-1:0] dout;							// 16 bits data [15:0] dout
 
 reg [DWIDTH-1:0] dout;                             //[15:0] dout sigmoid(addr)
 reg [DWIDTH_TMP-1:0] dout_tmp;	                    //[31:0] temporary signal for dout
 reg [DWIDTH_TMP-1:0] mem [0:(2**AWIDTH-1)];		// [31:0] mem [0:255]

 initial begin
			mem[8'b1000_0000]=32'b0000_0000_0000_0000_0001_0101_1111_1010;	//-8.0000
			mem[8'b1000_0001]=32'b0000_0000_0000_0000_0001_0111_0110_0101;
			mem[8'b1000_0010]=32'b0000_0000_0000_0000_0001_1000_1110_0111;
			mem[8'b1000_0011]=32'b0000_0000_0000_0000_0001_1010_1000_0010;
			mem[8'b1000_0100]=32'b0000_0000_0000_0000_0001_1100_0011_1000;
			mem[8'b1000_0101]=32'b0000_0000_0000_0000_0001_1110_0000_1001;
			mem[8'b1000_0110]=32'b0000_0000_0000_0000_0001_1111_1111_1001;
			mem[8'b1000_0111]=32'b0000_0000_0000_0000_0010_0010_0000_1000;
			mem[8'b1000_1000]=32'b0000_0000_0000_0000_0010_0100_0011_1010;
			mem[8'b1000_1001]=32'b0000_0000_0000_0000_0010_0110_1001_0000;
			mem[8'b1000_1010]=32'b0000_0000_0000_0000_0010_1001_0000_1100;
			mem[8'b1000_1011]=32'b0000_0000_0000_0000_0010_1011_1011_0001;
			mem[8'b1000_1100]=32'b0000_0000_0000_0000_0010_1110_1000_0010;
			mem[8'b1000_1101]=32'b0000_0000_0000_0000_0011_0001_1000_0010;
			mem[8'b1000_1110]=32'b0000_0000_0000_0000_0011_0100_1011_0010;
			mem[8'b1000_1111]=32'b0000_0000_0000_0000_0011_1000_0001_1000;
			//end at -7.06250
			mem[8'b1001_0000]=32'b0000_0000_0000_0000_0011_1011_1011_0101;	//-7.0000
			mem[8'b1001_0001]=32'b0000_0000_0000_0000_0011_1111_1000_1110;
			mem[8'b1001_0010]=32'b0000_0000_0000_0000_0100_0011_1010_0110;
			mem[8'b1001_0011]=32'b0000_0000_0000_0000_0100_1000_0000_0010;
			mem[8'b1001_0100]=32'b0000_0000_0000_0000_0100_1100_1010_0101;
			mem[8'b1001_0101]=32'b0000_0000_0000_0000_0101_0001_1001_0101;
			mem[8'b1001_0110]=32'b0000_0000_0000_0000_0101_0110_1101_0110;
			mem[8'b1001_0111]=32'b0000_0000_0000_0000_0101_1100_0110_0010;
			mem[8'b1001_1000]=32'b0000_0000_0000_0000_0110_0010_0110_0010;
			mem[8'b1001_1001]=32'b0000_0000_0000_0000_0110_1000_1011_0111;
			mem[8'b1001_1010]=32'b0000_0000_0000_0000_0110_1111_0111_0101;
			mem[8'b1001_1011]=32'b0000_0000_0000_0000_0111_0110_1010_0010;
			mem[8'b1001_1100]=32'b0000_0000_0000_0000_0111_1110_0100_0101;
			mem[8'b1001_1101]=32'b0000_0000_0000_0000_1000_0110_0110_0110;
			mem[8'b1001_1110]=32'b0000_0000_0000_0000_1000_1111_0000_1100;
			mem[8'b1001_1111]=32'b0000_0000_0000_0000_1001_1000_0100_0000;
			//end at -6.06250
			mem[8'b1010_0000]=32'b0000_0000_0000_0000_1010_0010_0000_1100;	//-6.0000
			mem[8'b1010_0001]=32'b0000_0000_0000_0000_1010_1100_0111_1000;
			mem[8'b1010_0010]=32'b0000_0000_0000_0000_1011_0111_1001_0000;
			mem[8'b1010_0011]=32'b0000_0000_0000_0000_1100_0011_0101_1101;
			mem[8'b1010_0100]=32'b0000_0000_0000_0000_1100_1111_1110_1101;
			mem[8'b1010_0101]=32'b0000_0000_0000_0000_1101_1101_0100_1010;
			mem[8'b1010_0110]=32'b0000_0000_0000_0000_1110_1011_1000_0011;
			mem[8'b1010_0111]=32'b0000_0000_0000_0000_1111_1010_1010_0100;
			mem[8'b1010_1000]=32'b0000_0000_0000_0001_0000_1010_1011_1110;
			mem[8'b1010_1001]=32'b0000_0000_0000_0001_0001_1011_1101_1111;
			mem[8'b1010_1010]=32'b0000_0000_0000_0001_0010_1110_0001_1000;
			mem[8'b1010_1011]=32'b0000_0000_0000_0001_0100_0001_0111_1011;
			mem[8'b1010_1100]=32'b0000_0000_0000_0001_0101_0110_0001_1011;
			mem[8'b1010_1101]=32'b0000_0000_0000_0001_0110_1100_0000_1100;
			mem[8'b1010_1110]=32'b0000_0000_0000_0001_1000_0011_0110_0011;
			mem[8'b1010_1111]=32'b0000_0000_0000_0001_1001_1100_0011_0111;
			//end at -5.06250
			mem[8'b1011_0000]=32'b0000_0000_0000_0001_1011_0110_1001_1111;	//-5.0000
			mem[8'b1011_0001]=32'b0000_0000_0000_0001_1101_0010_1011_0110;
			mem[8'b1011_0010]=32'b0000_0000_0000_0001_1111_0000_1001_0101;
			mem[8'b1011_0011]=32'b0000_0000_0000_0010_0001_0000_0101_1010;
			mem[8'b1011_0100]=32'b0000_0000_0000_0010_0011_0010_0010_0010;
			mem[8'b1011_0101]=32'b0000_0000_0000_0010_0101_0110_0000_1111;
			mem[8'b1011_0110]=32'b0000_0000_0000_0010_0111_1100_0100_0001;
			mem[8'b1011_0111]=32'b0000_0000_0000_0010_1010_0100_1101_1110;
			mem[8'b1011_1000]=32'b0000_0000_0000_0010_1101_0000_0000_1010;
			mem[8'b1011_1001]=32'b0000_0000_0000_0010_1111_1101_1111_0000;
			mem[8'b1011_1010]=32'b0000_0000_0000_0011_0010_1110_1011_1000;
			mem[8'b1011_1011]=32'b0000_0000_0000_0011_0110_0010_1001_0010;
			mem[8'b1011_1100]=32'b0000_0000_0000_0011_1001_1001_1010_1101;
			mem[8'b1011_1101]=32'b0000_0000_0000_0011_1101_0100_0011_1010;
			mem[8'b1011_1110]=32'b0000_0000_0000_0100_0001_0010_0111_0001;
			mem[8'b1011_1111]=32'b0000_0000_0000_0100_0101_0100_1000_1001;
			//end at -4.06250
			mem[8'b1100_0000]=32'b0000_0000_0000_0100_1001_1010_1011_1111;	//-4.0000
			mem[8'b1100_0001]=32'b0000_0000_0000_0100_1110_0101_0101_0000;
			mem[8'b1100_0010]=32'b0000_0000_0000_0101_0011_0100_1000_0000;
			mem[8'b1100_0011]=32'b0000_0000_0000_0101_1000_1000_1001_0101;
			mem[8'b1100_0100]=32'b0000_0000_0000_0101_1110_0001_1101_1000;
			mem[8'b1100_0101]=32'b0000_0000_0000_0110_0100_0000_1001_0111;
			mem[8'b1100_0110]=32'b0000_0000_0000_0110_1010_0101_0010_0100;
			mem[8'b1100_0111]=32'b0000_0000_0000_0111_0000_1111_1101_0100;
			mem[8'b1100_1000]=32'b0000_0000_0000_0111_1000_0001_0000_0010;
			mem[8'b1100_1001]=32'b0000_0000_0000_0111_1111_1001_0000_0011;
			mem[8'b1100_1010]=32'b0000_0000_0000_1000_0111_1000_0100_0011;
			mem[8'b1100_1011]=32'b0000_0000_0000_1000_1111_1111_0100_0001;
			mem[8'b1100_1100]=32'b0000_0000_0000_1001_1000_1110_0100_0001;
			mem[8'b1100_1101]=32'b0000_0000_0000_1010_0010_0101_1100_0101;
			mem[8'b1100_1110]=32'b0000_0000_0000_1010_1100_0110_0100_0011;
			mem[8'b1100_1111]=32'b0000_0000_0000_1011_0111_0000_0011_0101;
			//end at -3.06250
			mem[8'b1101_0000]=32'b0000_0000_0000_1100_0010_0100_0001_1010;	//-3.0000
			mem[8'b1101_0001]=32'b0000_0000_0000_1100_1110_0010_0111_1000;
			mem[8'b1101_0010]=32'b0000_0000_0000_1101_1010_1011_1101_0111;
			mem[8'b1101_0011]=32'b0000_0000_0000_1110_1000_0000_1100_0110;
			mem[8'b1101_0100]=32'b0000_0000_0000_1111_0110_0001_1101_0111;
			mem[8'b1101_0101]=32'b0000_0000_0001_0000_0100_1111_1010_0000;
			mem[8'b1101_0110]=32'b0000_0000_0001_0001_0100_1010_1011_1101;
			mem[8'b1101_0111]=32'b0000_0000_0001_0010_0101_0011_1100_1101;
			mem[8'b1101_1000]=32'b0000_0000_0001_0011_0110_1011_0111_0001;
			mem[8'b1101_1001]=32'b0000_0000_0001_0100_1001_0010_0100_1111;
			mem[8'b1101_1010]=32'b0000_0000_0001_0101_1100_1001_0000_1101;
			mem[8'b1101_1011]=32'b0000_0000_0001_0111_0001_0000_0101_0110;
			mem[8'b1101_1100]=32'b0000_0000_0001_1000_0110_1000_1101_0011;
			mem[8'b1101_1101]=32'b0000_0000_0001_1001_1101_0011_0010_1110;
			mem[8'b1101_1110]=32'b0000_0000_0001_1011_0101_0000_0001_0011;
			mem[8'b1101_1111]=32'b0000_0000_0001_1100_1110_0000_0010_1001;
			//end at -2.06250
			mem[8'b1110_0000]=32'b00000000000111101000010000010101;	//-2.0000
			mem[8'b1110_0001]=32'b00000000001000000011110001111001;
			mem[8'b1110_0010]=32'b00000000001000100000100111110010;
			mem[8'b1110_0011]=32'b00000000001000111110110100010100;
			mem[8'b1110_0100]=32'b00000000001001011110011001101100;
			mem[8'b1110_0101]=32'b00000000001001111111011001111110;
			mem[8'b1110_0110]=32'b00000000001010100001110111000000;
			mem[8'b1110_0111]=32'b00000000001011000101110010011110;
			mem[8'b1110_1000]=32'b00000000001011101011001101110000;
			mem[8'b1110_1001]=32'b00000000001100010010001010000010;
			mem[8'b1110_1010]=32'b00000000001100111010101000001000;
			mem[8'b1110_1011]=32'b00000000001101100100101000100100;
			mem[8'b1110_1100]=32'b00000000001110010000001011100000;
			mem[8'b1110_1101]=32'b00000000001110111101010000101110;
			mem[8'b1110_1110]=32'b00000000001111101011110111100100;
			mem[8'b1110_1111]=32'b00000000010000011011111110111110;
			//end at -1.06250
			mem[8'b1111_0000]=32'b00000000010001001101100101011000;	//-1.0000
			mem[8'b1111_0001]=32'b00000000010010000000101000110011;
			mem[8'b1111_0010]=32'b00000000010010110101000110101100;
			mem[8'b1111_0011]=32'b00000000010011101010111100000100;
			mem[8'b1111_0100]=32'b00000000010100100010000101011000;
			mem[8'b1111_0101]=32'b00000000010101011010011110100111;
			mem[8'b1111_0110]=32'b00000000010110010100000011001111;
			mem[8'b1111_0111]=32'b00000000010111001110101110001101;
			mem[8'b1111_1000]=32'b00000000011000001010011010000001;
			mem[8'b1111_1001]=32'b00000000011001000111000000110000;
			mem[8'b1111_1010]=32'b00000000011010000100011100000000;
			mem[8'b1111_1011]=32'b00000000011011000010100101000100;
			mem[8'b1111_1100]=32'b00000000011100000001010100110011;
			mem[8'b1111_1101]=32'b00000000011101000000100011111000;
			mem[8'b1111_1110]=32'b00000000011110000000001010101010;
			mem[8'b1111_1111]=32'b00000000011111000000000001010101;
			//end at -0.06250
			mem[8'b0000_0000]=32'b00000000100000000000000000000000;	//0.0000
			mem[8'b0000_0001]=32'b00000000100000111111111110101011;
			mem[8'b0000_0010]=32'b00000000100001111111110101010110;
			mem[8'b0000_0011]=32'b00000000100010111111011100001000;
			mem[8'b0000_0100]=32'b00000000100011111110101011001101;
			mem[8'b0000_0101]=32'b00000000100100111101011010111100;
			mem[8'b0000_0110]=32'b00000000100101111011100100000000;
			mem[8'b0000_0111]=32'b00000000100110111000111111010000;
			mem[8'b0000_1000]=32'b00000000100111110101100101111111;
			mem[8'b0000_1001]=32'b00000000101000110001010001110011;
			mem[8'b0000_1010]=32'b00000000101001101011111100110001;
			mem[8'b0000_1011]=32'b00000000101010100101100001011001;
			mem[8'b0000_1100]=32'b00000000101011011101111010101000;
			mem[8'b0000_1101]=32'b00000000101100010101000011111100;
			mem[8'b0000_1110]=32'b00000000101101001010111001010100;
			mem[8'b0000_1111]=32'b00000000101101111111010111001101;
			//end at 0.93750
			mem[8'b0001_0000]=32'b00000000101110110010011010101000;	//1.0000
			mem[8'b0001_0001]=32'b00000000101111100100000001000010;
			mem[8'b0001_0010]=32'b00000000110000010100001000011100;
			mem[8'b0001_0011]=32'b00000000110001000010101111010010;
			mem[8'b0001_0100]=32'b00000000110001101111110100100000;
			mem[8'b0001_0101]=32'b00000000110010011011010111011100;
			mem[8'b0001_0110]=32'b00000000110011000101010111111000;
			mem[8'b0001_0111]=32'b00000000110011101101110101111110;
			mem[8'b0001_1000]=32'b00000000110100010100110010010000;
			mem[8'b0001_1001]=32'b00000000110100111010001101100010;
			mem[8'b0001_1010]=32'b00000000110101011110001001000000;
			mem[8'b0001_1011]=32'b00000000110110000000100110000010;
			mem[8'b0001_1100]=32'b00000000110110100001100110010100;
			mem[8'b0001_1101]=32'b00000000110111000001001011101100;
			mem[8'b0001_1110]=32'b00000000110111011111011000001110;
			mem[8'b0001_1111]=32'b00000000110111111100001110000111;
			//end at 1.93750
			mem[8'b0010_0000]=32'b00000000111000010111101111101011;	//2.0000
			mem[8'b0010_0001]=32'b00000000111000110001111111010111;
			mem[8'b0010_0010]=32'b00000000111001001010111111101101;
			mem[8'b0010_0011]=32'b00000000111001100010110011010010;
			mem[8'b0010_0100]=32'b00000000111001111001011100101101;
			mem[8'b0010_0101]=32'b00000000111010001110111110101010;
			mem[8'b0010_0110]=32'b00000000111010100011011011110011;
			mem[8'b0010_0111]=32'b00000000111010110110110110110001;
			mem[8'b0010_1000]=32'b00000000111011001001010010001111;
			mem[8'b0010_1001]=32'b00000000111011011010110000110011;
			mem[8'b0010_1010]=32'b00000000111011101011010101000011;
			mem[8'b0010_1011]=32'b00000000111011111011000001100000;
			mem[8'b0010_1100]=32'b00000000111100001001111000101001;
			mem[8'b0010_1101]=32'b00000000111100010111111100111010;
			mem[8'b0010_1110]=32'b00000000111100100101010000101001;
			mem[8'b0010_1111]=32'b00000000111100110001110110001000;
			//end at 2.93750
			mem[8'b0011_0000]=32'b00000000111100111101101111100110;	//3.0000
			mem[8'b0011_0001]=32'b00000000111101001000111111001011;
			mem[8'b0011_0010]=32'b00000000111101010011100110111101;
			mem[8'b0011_0011]=32'b00000000111101011101101000111011;
			mem[8'b0011_0100]=32'b00000000111101100111000110111111;
			mem[8'b0011_0101]=32'b00000000111101110000000010111111;
			mem[8'b0011_0110]=32'b00000000111101111000011110101101;
			mem[8'b0011_0111]=32'b00000000111110000000011011110101;
			mem[8'b0011_1000]=32'b00000000111110000111111011111110;
			mem[8'b0011_1001]=32'b00000000111110001111000000101100;
			mem[8'b0011_1010]=32'b00000000111110010101101011011100;
			mem[8'b0011_1011]=32'b00000000111110011011111101101001;
			mem[8'b0011_1100]=32'b00000000111110100001111000101000;
			mem[8'b0011_1101]=32'b00000000111110100111011101101011;
			mem[8'b0011_1110]=32'b00000000111110101100101110000000;
			mem[8'b0011_1111]=32'b00000000111110110001101010110000;
			//end at 3.93750
			mem[8'b0100_0000]=32'b00000000111110110110010101000001;	//4.0000
			mem[8'b0100_0001]=32'b00000000111110111010101101110111;
			mem[8'b0100_0010]=32'b00000000111110111110110110001111;
			mem[8'b0100_0011]=32'b00000000111111000010101111000110;
			mem[8'b0100_0100]=32'b00000000111111000110011001010011;
			mem[8'b0100_0101]=32'b00000000111111001001110101101110;
			mem[8'b0100_0110]=32'b00000000111111001101000101001000;
			mem[8'b0100_0111]=32'b00000000111111010000001000010000;
			mem[8'b0100_1000]=32'b00000000111111010010111111110110;
			mem[8'b0100_1001]=32'b00000000111111010101101100100010;
			mem[8'b0100_1010]=32'b00000000111111011000001110111111;
			mem[8'b0100_1011]=32'b00000000111111011010100111110001;
			mem[8'b0100_1100]=32'b00000000111111011100110111011110;
			mem[8'b0100_1101]=32'b00000000111111011100110111011110;
			mem[8'b0100_1110]=32'b00000000111111100000111101101011;
			mem[8'b0100_1111]=32'b00000000111111100010110101001010;
			//end at 4.93750
			mem[8'b0101_0000]=32'b00000000111111100100100101100001;	//5.0000
			mem[8'b0101_0001]=32'b00000000111111100110001111001001;
			mem[8'b0101_0010]=32'b00000000111111100111110010011101;
			mem[8'b0101_0011]=32'b00000000111111101001001111110100;
			mem[8'b0101_0100]=32'b00000000111111101010100111100101;
			mem[8'b0101_0101]=32'b00000000111111101011111010000101;
			mem[8'b0101_0110]=32'b00000000111111101101000111101000;
			mem[8'b0101_0111]=32'b00000000111111101110010000100001;
			mem[8'b0101_1000]=32'b00000000111111101111010101000010;
			mem[8'b0101_1001]=32'b00000000111111110000010101011100;
			mem[8'b0101_1010]=32'b00000000111111110001010001111101;
			mem[8'b0101_1011]=32'b00000000111111110010001010110110;
			mem[8'b0101_1100]=32'b00000000111111110011000000010011;
			mem[8'b0101_1101]=32'b00000000111111110011110010100011;
			mem[8'b0101_1110]=32'b00000000111111110100100001110000;
			mem[8'b0101_1111]=32'b00000000111111110101001110001000;
			//end at 5.93750
			mem[8'b0110_0000]=32'b00000000111111110101110111110100;	//6.0000
			mem[8'b0110_0001]=32'b00000000111111110110011111000000;
			mem[8'b0110_0010]=32'b00000000111111110111000011110100;
			mem[8'b0110_0011]=32'b00000000111111110111100110011010;
			mem[8'b0110_0100]=32'b00000000111111111000000110111011;
			mem[8'b0110_0101]=32'b00000000111111111000100101011110;
			mem[8'b0110_0110]=32'b00000000111111111001000010001011;
			mem[8'b0110_0111]=32'b00000000111111111001011101001001;
			mem[8'b0110_1000]=32'b00000000111111111001110110011110;
			mem[8'b0110_1001]=32'b00000000111111111010001110010010;
			mem[8'b0110_1010]=32'b00000000111111111010100100101010;
			mem[8'b0110_1011]=32'b00000000111111111010111001101011;
			mem[8'b0110_1100]=32'b00000000111111111011001101011011;
			mem[8'b0110_1101]=32'b00000000111111111011011111111110;
			mem[8'b0110_1110]=32'b00000000111111111011110001011010;
			mem[8'b0110_1111]=32'b00000000111111111100000001110010;
			//end at 6.93750
			mem[8'b0111_0000]=32'b00000000111111111100010001001011;	//7.0000
			mem[8'b0111_0001]=32'b00000000111111111100011111101000;
			mem[8'b0111_0010]=32'b00000000111111111100101101001110;
			mem[8'b0111_0011]=32'b00000000111111111100111001111110;
			mem[8'b0111_0100]=32'b00000000111111111101000101111110;
			mem[8'b0111_0101]=32'b00000000111111111101010001001111;
			mem[8'b0111_0110]=32'b00000000111111111101011011110100;
			mem[8'b0111_0111]=32'b00000000111111111101100101110000;
			mem[8'b0111_1000]=32'b00000000111111111101101111000110;
			mem[8'b0111_1001]=32'b00000000111111111101110111111000;
			mem[8'b0111_1010]=32'b00000000111111111110000000000111;
			mem[8'b0111_1011]=32'b00000000111111111110000111110111;
			mem[8'b0111_1100]=32'b00000000111111111110001111001000;
			mem[8'b0111_1101]=32'b00000000111111111110010101111110;
			mem[8'b0111_1110]=32'b00000000111111111110011100011001;
			mem[8'b0111_1111]=32'b00000000111111111110100010011011;
			//end at 7.93750
end
 
 always@(posedge clk) begin
   if(din==1) 						//only READ is used
	begin
		dout_tmp = mem[addr]; 	    //0000_0000.0000_0000_0000_0000_0000_0000
		dout = dout_tmp[29:14];	    //00_0000.0000_0000_00
	end
	else 
		dout = 16'bz;				//when no control signal is given, tristate the output
	end

endmodule
 
