-------------------------------------------------------------------------------
-- Title      : Linear feedback shift register
-- Project    : 
-------------------------------------------------------------------------------
-- File       : lfsr.vhd
-- Author     : Hieu D. Bui  <Hieu D. Bui@>
-- Company    : SISLAB, VNU-UET
-- Created    : 2017-12-14
-- Last update: 2017-12-15
-- Platform   : 
-- Standard   : VHDL'08
-------------------------------------------------------------------------------
-- Description: A generic linear feedback ship register for stochastic
--              computing
-------------------------------------------------------------------------------
-- Copyright (c) 2017 SISLAB, VNU-UET
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2017-12-14  1.0      Hieu D. Bui     Created
-------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY lfsr IS

  GENERIC (
    DATA_WIDTH : INTEGER := 8);

  PORT (
    clk         : IN  STD_LOGIC;
    rst_n       : IN  STD_LOGIC;
    seed_in     : IN  STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
    set_seed_in : IN  STD_LOGIC;
    enable_in   : IN  STD_LOGIC;
    lfsr_out    : OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));

END ENTITY lfsr;


ARCHITECTURE beh OF lfsr IS
  TYPE int_array_t IS ARRAY (0 TO 6) OF INTEGER;
  TYPE int_array_2d_t IS ARRAY (NATURAL RANGE <>) OF int_array_t;
  -- the following constants are taken from
  -- https://www.xilinx.com/support/documentation/application_notes/xapp052.pdf
  -- this file implement maximum length lfsr using xnor function
  -- content of the lfsr should not be all '1's
  -- the index of the array is the number of bits of the lfsr
  -- the first index of the subarray: number of taps
  -- the following indexs of the subarray: taps' posistions
  -- 0 indicates that the index is not used
  CONSTANT lfsr_taps : int_array_2d_t(3 TO 168)
    -- numTaps
    := (
      (2, 3, 2, 0, 0, 0, 0),            -- 3
      (2, 4, 3, 0, 0, 0, 0),            -- 4
      (2, 5, 3, 0, 0, 0, 0),            -- 5
      (2, 6, 5, 0, 0, 0, 0),            -- 6
      (2, 7, 6, 0, 0, 0, 0),            -- 7
      (4, 8, 6, 5, 4, 0, 0),            -- 8
      (2, 9, 5, 0, 0, 0, 0),            -- 9
      (2, 10, 7, 0, 0, 0, 0),           -- 10
      (2, 11, 9, 0, 0, 0, 0),           -- 11
      (4, 12, 6, 4, 1, 0, 0),           -- 12
      (4, 13, 4, 3, 1, 0, 0),           -- 13
      (4, 14, 5, 3, 1, 0, 0),           -- 14
      (2, 15, 14, 0, 0, 0, 0),          -- 15
      (4, 16, 15, 13, 4, 0, 0),         -- 16
      (2, 17, 14, 0, 0, 0, 0),          -- 17
      (2, 18, 11, 0, 0, 0, 0),          -- 18
      (4, 19, 6, 2, 1, 0, 0),           -- 19
      (2, 20, 17, 0, 0, 0, 0),          -- 20
      (2, 21, 19, 0, 0, 0, 0),          -- 21
      (2, 22, 21, 0, 0, 0, 0),          -- 22
      (2, 23, 18, 0, 0, 0, 0),          -- 23
      (4, 24, 23, 22, 17, 0, 0),        -- 24
      (2, 25, 22, 0, 0, 0, 0),          -- 25
      (4, 26, 6, 2, 1, 0, 0),           -- 26
      (4, 27, 5, 2, 1, 0, 0),           -- 27
      (2, 28, 25, 0, 0, 0, 0),          -- 28
      (2, 29, 27, 0, 0, 0, 0),          -- 29
      (4, 30, 6, 4, 1, 0, 0),           -- 30
      (2, 31, 28, 0, 0, 0, 0),          -- 31
      (4, 32, 22, 2, 1, 0, 0),          -- 32
      (2, 33, 20, 0, 0, 0, 0),          -- 33
      (4, 34, 27, 2, 1, 0, 0),          -- 34
      (2, 35, 33, 0, 0, 0, 0),          -- 35
      (2, 36, 25, 0, 0, 0, 0),          -- 36
      (6, 37, 5, 4, 3, 2, 1),           -- 37
      (4, 38, 6, 5, 1, 0, 0),           -- 38
      (2, 39, 35, 0, 0, 0, 0),          -- 39
      (4, 40, 38, 21, 19, 0, 0),        -- 40
      (2, 41, 38, 0, 0, 0, 0),          -- 41
      (4, 42, 41, 20, 19, 0, 0),        -- 42
      (4, 43, 42, 38, 37, 0, 0),        -- 43
      (4, 44, 43, 18, 17, 0, 0),        -- 44
      (4, 45, 44, 42, 41, 0, 0),        -- 45
      (4, 46, 45, 26, 25, 0, 0),        -- 46
      (2, 47, 42, 0, 0, 0, 0),          -- 47
      (4, 48, 47, 21, 20, 0, 0),        -- 48
      (2, 49, 40, 0, 0, 0, 0),          -- 49
      (4, 50, 49, 24, 23, 0, 0),        -- 50
      (4, 51, 50, 36, 35, 0, 0),        -- 51
      (2, 52, 49, 0, 0, 0, 0),          -- 52
      (4, 53, 52, 38, 37, 0, 0),        -- 53
      (4, 54, 53, 18, 17, 0, 0),        -- 54
      (2, 55, 31, 0, 0, 0, 0),          -- 55
      (4, 56, 55, 35, 34, 0, 0),        -- 56
      (2, 57, 50, 0, 0, 0, 0),          -- 57
      (2, 58, 39, 0, 0, 0, 0),          -- 58
      (4, 59, 58, 38, 37, 0, 0),        -- 59
      (2, 60, 59, 0, 0, 0, 0),          -- 60
      (4, 61, 60, 46, 45, 0, 0),        -- 61
      (4, 62, 61, 6, 5, 0, 0),          -- 62
      (2, 63, 62, 0, 0, 0, 0),          -- 63
      (4, 64, 63, 61, 60, 0, 0),        -- 64
      (2, 65, 47, 0, 0, 0, 0),          -- 65
      (4, 66, 65, 57, 56, 0, 0),        -- 66
      (4, 67, 66, 58, 57, 0, 0),        -- 67
      (2, 68, 59, 0, 0, 0, 0),          -- 68
      (4, 69, 67, 42, 40, 0, 0),        -- 69
      (4, 70, 69, 55, 54, 0, 0),        -- 70
      (2, 71, 65, 0, 0, 0, 0),          -- 71
      (4, 72, 66, 25, 19, 0, 0),        -- 72
      (2, 73, 48, 0, 0, 0, 0),          -- 73
      (4, 74, 73, 59, 58, 0, 0),        -- 74
      (4, 75, 74, 65, 64, 0, 0),        -- 75
      (4, 76, 75, 41, 40, 0, 0),        -- 76
      (4, 77, 76, 47, 46, 0, 0),        -- 77
      (4, 78, 77, 59, 58, 0, 0),        -- 78
      (2, 79, 70, 0, 0, 0, 0),          -- 79
      (4, 80, 79, 43, 42, 0, 0),        -- 80
      (2, 81, 77, 0, 0, 0, 0),          -- 81
      (4, 82, 79, 47, 44, 0, 0),        -- 82
      (4, 83, 82, 38, 37, 0, 0),        -- 83
      (2, 84, 71, 0, 0, 0, 0),          -- 84
      (4, 85, 84, 58, 57, 0, 0),        -- 85
      (4, 86, 85, 74, 73, 0, 0),        -- 86
      (2, 87, 74, 0, 0, 0, 0),          -- 87
      (4, 88, 87, 17, 16, 0, 0),        -- 88
      (2, 89, 51, 0, 0, 0, 0),          -- 89
      (4, 90, 89, 72, 71, 0, 0),        -- 90
      (4, 91, 90, 8, 7, 0, 0),          -- 91
      (4, 92, 91, 80, 79, 0, 0),        -- 92
      (2, 93, 91, 0, 0, 0, 0),          -- 93
      (2, 94, 73, 0, 0, 0, 0),          -- 94
      (2, 95, 84, 0, 0, 0, 0),          -- 95
      (4, 96, 94, 49, 47, 0, 0),        -- 96
      (2, 97, 91, 0, 0, 0, 0),          -- 97
      (2, 98, 87, 0, 0, 0, 0),          -- 98
      (4, 99, 97, 54, 52, 0, 0),        -- 99
      (2, 100, 63, 0, 0, 0, 0),         -- 100
      (4, 101, 100, 95, 94, 0, 0),      -- 101
      (4, 102, 101, 36, 35, 0, 0),      -- 102
      (2, 103, 94, 0, 0, 0, 0),         -- 103
      (4, 104, 103, 94, 93, 0, 0),      -- 104
      (2, 105, 89, 0, 0, 0, 0),         -- 105
      (2, 106, 91, 0, 0, 0, 0),         -- 106
      (4, 107, 105, 44, 42, 0, 0),      -- 107
      (2, 108, 77, 0, 0, 0, 0),         -- 108
      (4, 109, 108, 103, 102, 0, 0),    -- 109
      (4, 110, 109, 98, 97, 0, 0),      -- 110
      (2, 111, 101, 0, 0, 0, 0),        -- 111
      (4, 112, 110, 69, 67, 0, 0),      -- 112
      (2, 113, 104, 0, 0, 0, 0),        -- 113
      (4, 114, 113, 33, 32, 0, 0),      -- 114
      (4, 115, 114, 101, 100, 0, 0),    -- 115
      (4, 116, 115, 46, 45, 0, 0),      -- 116
      (4, 117, 115, 99, 97, 0, 0),      -- 117
      (2, 118, 85, 0, 0, 0, 0),         -- 118
      (2, 119, 111, 0, 0, 0, 0),        -- 119
      (4, 120, 113, 9, 2, 0, 0),        -- 120
      (2, 121, 103, 0, 0, 0, 0),        -- 121
      (4, 122, 121, 63, 62, 0, 0),      -- 122
      (2, 123, 121, 0, 0, 0, 0),        -- 123
      (2, 124, 87, 0, 0, 0, 0),         -- 124
      (4, 125, 124, 18, 17, 0, 0),      -- 125
      (4, 126, 125, 90, 89, 0, 0),      -- 126
      (2, 127, 126, 0, 0, 0, 0),        -- 127
      (4, 128, 126, 101, 99, 0, 0),     -- 128
      (2, 129, 124, 0, 0, 0, 0),        -- 129
      (2, 130, 127, 0, 0, 0, 0),        -- 130
      (4, 131, 130, 84, 83, 0, 0),      -- 131
      (2, 132, 103, 0, 0, 0, 0),        -- 132
      (4, 133, 132, 82, 81, 0, 0),      -- 133
      (2, 134, 77, 0, 0, 0, 0),         -- 134
      (2, 135, 124, 0, 0, 0, 0),        -- 135
      (4, 136, 135, 11, 10, 0, 0),      -- 136
      (2, 137, 116, 0, 0, 0, 0),        -- 137
      (4, 138, 137, 131, 130, 0, 0),    -- 138
      (4, 139, 136, 134, 131, 0, 0),    -- 139
      (2, 140, 111, 0, 0, 0, 0),        -- 140
      (4, 141, 140, 110, 109, 0, 0),    -- 141
      (2, 142, 121, 0, 0, 0, 0),        -- 142
      (4, 143, 142, 123, 122, 0, 0),    -- 143
      (4, 144, 143, 75, 74, 0, 0),      -- 144
      (2, 145, 93, 0, 0, 0, 0),         -- 145
      (4, 146, 145, 87, 86, 0, 0),      -- 146
      (4, 147, 146, 110, 109, 0, 0),    -- 147
      (2, 148, 121, 0, 0, 0, 0),        -- 148
      (4, 149, 148, 40, 39, 0, 0),      -- 149
      (2, 150, 97, 0, 0, 0, 0),         -- 150
      (2, 151, 148, 0, 0, 0, 0),        -- 151
      (4, 152, 151, 87, 86, 0, 0),      -- 152
      (2, 153, 152, 0, 0, 0, 0),        -- 153
      (4, 154, 152, 27, 25, 0, 0),      -- 154
      (4, 155, 154, 124, 123, 0, 0),    -- 155
      (4, 156, 155, 41, 40, 0, 0),      -- 156
      (4, 157, 156, 131, 130, 0, 0),    -- 157
      (4, 158, 157, 132, 131, 0, 0),    -- 158
      (2, 159, 128, 0, 0, 0, 0),        -- 159
      (4, 160, 159, 142, 141, 0, 0),    -- 160
      (2, 161, 143, 0, 0, 0, 0),        -- 161
      (4, 162, 161, 75, 74, 0, 0),      -- 162
      (4, 163, 162, 104, 103, 0, 0),    -- 163
      (4, 164, 163, 151, 150, 0, 0),    -- 164
      (4, 165, 164, 135, 134, 0, 0),    -- 165
      (4, 166, 165, 128, 127, 0, 0),    -- 166
      (2, 167, 161, 0, 0, 0, 0),        -- 167
      (4, 168, 166, 153, 151, 0, 0)     -- 168
      );
  SIGNAL lfsr_reg        : STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL lfsr_feedback   : STD_LOGIC;
  SIGNAL feedback_vector : STD_LOGIC_VECTOR(lfsr_taps(DATA_WIDTH)(0)-1 DOWNTO 0);
BEGIN  -- ARCHITECTURE beh

  feedback_gen : FOR i IN 0 TO lfsr_taps(DATA_WIDTH)(0)-1 GENERATE
    feedback_vector(i) <= lfsr_reg(lfsr_taps(DATA_WIDTH)(i+1)-1);
  END GENERATE feedback_gen;

  lfsr_feedback <= XNOR(feedback_vector);

  lfsr_proc : PROCESS (clk, rst_n) IS
  BEGIN  -- PROCESS lfsr_proc
    IF rst_n = '0' THEN                 -- asynchronous reset (active low)
      lfsr_reg <= (OTHERS => '0');
    ELSIF rising_edge(clk) THEN         -- rising clock edge
      IF set_seed_in = '1' THEN
        lfsr_reg <= seed_in;
        --pragma synthesis_off
        ASSERT nand(seed_in) REPORT "Illegal seed value" SEVERITY FAILURE;
        --pragma synthesis_on
      ELSIF enable_in = '1' THEN
        lfsr_reg <= lfsr_reg(DATA_WIDTH-2 DOWNTO 0) & lfsr_feedback;
      END IF;
    END IF;
  END PROCESS lfsr_proc;

  lfsr_out <= lfsr_reg;
END ARCHITECTURE beh;
